library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity channel is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity channel;

architecture RTL of channel is
    
begin

end architecture RTL;
