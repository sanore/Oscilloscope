library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity channel_tb is
end entity channel_tb;

architecture RTL of channel_tb is
    
begin

end architecture RTL;
