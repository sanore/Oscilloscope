library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity ram;

architecture RTL of ram is
    
begin

end architecture RTL;
