library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrlunit_tb_tb is
end entity ctrlunit_tb_tb;

architecture RTL of ctrlunit_tb_tb is
component ctrlunit
    generic(
        ADDR_WIDTH : integer := 13;
        DATA_WIDTH : integer := 16
    );
    port(
        clk           : in  std_logic;
        rst           : in  std_logic;
        start_record  : in  std_logic;
        adc_val       : in  std_ulogic_vector(11 downto 0);
        trigger_pulse : in  std_ulogic;
        write_address : out std_ulogic_vector(ADDR_WIDTH - 1 downto 0);
        write_data    : out std_ulogic_vector(DATA_WIDTH - 1 downto 0);
        write_en      : out std_ulogic;
        trigger_index : out std_ulogic_vector(ADDR_WIDTH - 1 downto 0)
    );
end component ctrlunit;
signal clk     : std_logic := '0';
signal reset   : std_logic := '1';
signal start   : std_logic := '0';
signal dut_adc_val : std_ulogic_vector(11 downto 0);
signal dut_trigger_pulse : std_ulogic := '0';

signal dut_write_address : std_ulogic_vector(13 - 1 downto 0);
signal dut_write_data    : std_ulogic_vector(16 - 1 downto 0);
signal dut_write_en      : std_ulogic;
signal dut_trigger_index : std_ulogic_vector(16 - 1 downto 0);
begin
    clk <= clk after 5 ns;
    reset <= '1', '0' after 50 ns;
    start <= '0', '1' after 100 ns;
    dut_trigger_pulse <= '0', '1' after 2 us, '0' after 10 ns;
dut:component ctrlunit
    port map(
        clk           => clk,
        rst           => reset,
        start_record  => start,
        adc_val       => dut_adc_val,
        trigger_pulse => dut_trigger_pulse,
        write_address => dut_write_address,
        write_data    => dut_write_data,
        write_en      => dut_write_en,
        trigger_index => dut_trigger_index
    ) ;
dut_state : process is
begin
    wait for 10 ns;
    assert(dut_write_en = '0');
    assert(dut_write_address = "000000000000");
    assert(dut_write_data = "0000000000000000");
    wait for 105 ns;
    assert(dut_write_en = '1');
    wait for 1 us;
    assert(dut_write_address = "0000000000001");
    wait for 2 us + 10 ns;
    assert dut_write_address = dut_trigger_index report "dut_trigger_index wrong" severity error;
    wait for 1 us;
    assert(dut_write_address = std_ulogic_vector(unsigned(dut_trigger_index) + 1));
end process dut_state;

end architecture RTL;
