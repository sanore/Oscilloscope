library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity trigger is
    port(
        clk           : in std_logic;
        rst           : in std_logic
    );
end entity trigger;

architecture RTL of trigger is

begin

end architecture RTL;
