library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity trigger_tb is
end entity trigger_tb;

architecture RTL of trigger_tb is
    
begin

end architecture RTL;
