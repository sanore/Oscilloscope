library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity osci is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity osci;

architecture RTL of osci is
    
begin

end architecture RTL;
