library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity osci_tb is
end entity osci_tb;

architecture RTL of osci_tb is
    
begin

end architecture RTL;
