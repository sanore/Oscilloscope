library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrlunit is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity ctrlunit;

architecture RTL of ctrlunit is
    
begin

end architecture RTL;
